* DC analysis on a simple circuit network

v1 a 0 dc 9
r1 a 0 5k
.op
.end
