* L08_P13 PoC
* plot -l(A)

r1 0 A 0.5k
l1 A 0 10m ic = 10m

.tran 10u 100u uic
.end
