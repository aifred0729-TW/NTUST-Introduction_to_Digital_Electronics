* L07_P17 PoC
* plot c(A)

r1 0 A 1k
c1 A 0 100u ic = 100u

.tran 10m 100m uic
.end
